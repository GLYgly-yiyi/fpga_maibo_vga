`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/11/14 18:17:33
// Design Name: 
// Module Name: rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module rom(
input wire[7:0] addr,
output wire[0:127] M
    );
    reg[0:127] rom[0:255];
    
    parameter data={
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111,//1
    
    
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100,//1
    
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000,//1
    
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000,//1
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000,//1
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000,//1
    
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000,//1
    
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000,//1
    
    
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000,//1
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000,//1
    
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000,//1
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000,//1
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000,//1
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000,//1
    
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000,//1
    
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000,//1
    
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000,//1
    
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000,//1
    
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000,//1
    
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000,//1
    
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000,//1
    
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000,//1
    
    
    128'b00000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    
    128'b00000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    
    128'b00000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    
    128'b00000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    
    128'b00000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    
    128'b00000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    128'b00111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b00111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b01110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b01110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    
    
    
    128'b11100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b11100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b11100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,//1
    128'b11100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000//1
    
    };
    integer i;
    initial
     begin
    for(i=0;i<256;i=i+1)
      rom[i]=data[(32767-128*i)-:128];
    end
    
    assign M=rom[addr];

    
    
endmodule
