`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/11/17 13:53:52
// Design Name: 
// Module Name: Fre_Vopp_mapping_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Fre_Vopp_mapping_rom(
   input wire[5:0]addr_Fre_Vopp,
output wire[0:63]F
    );
    
   reg[0:63]rom[0:63];
    
    parameter data={
    64'b0000000111111111111111000000000000000000000000000000000000000000,
    64'b0000000111111111111111000000000000000000000000000000000000000000,
    64'b0000000111000000000000000000000000000000000000000000000000000000,
    64'b0000000111000000000000000000000000000000000000000000000000000000,
    64'b0000000111000000000000000000000000000000000000000000000000000000,
    64'b0000000111000000000000000000000000000000000000000000000000000000,
    64'b0000000111000000000000000000000000000000000000000000000000000000,
    64'b0000000111000000000000000000000000000000000000000000000000000000,//7
    64'b0000000111000000000000000000000000000000000000000000000000000000,
    64'b0000000111000000000000000000000000000000000000000000000000000000,//9
    64'b0000000111000000000000000000000000000000000000000000000000000000,
    64'b0000000111000000000000000000000000000000000000000000000000000000,
    64'b0000000111000000000000000000000000000000000000000000000000000000,
    64'b0000000111000000000000000000000000000000000000000000000000000000,
    64'b0000000111000000000000000000000000000000000000000000000000000000,
    64'b0000000111111111111111000000000000000000000000000000000000000000,
    
    64'b0000000111111111111111000000010010000000010111111111101000001111,
    64'b0000000111000000000000000000010010000000010000000000101000001111,
    64'b0000000111000000000000000000100010000000010000000001000100001111,
    64'b0000000111000000000000000000100010000000010000000010000100001111,
    64'b0000000111000000000000000001000010000000010000000100000010000000,
    64'b0000000111000000000000000001000010000000010000000100000010000000,
    64'b0000000111000000000000000001000010000000010000001000000010000000,
    64'b0000000111000000000000000001000011111111110000010000000010000000,//7
    64'b0000000111000000000000000001000010000000010000010000000010000000,
    64'b0000000111000000000000000001000010000000010000100000000010000000,//9
    64'b0000000111000000000000000001000010000000010000100000000010000000,
    64'b0000000111000000000000000001000010000000010001000000000010000000,
    64'b0000000111000000000000000000100010000000010001000000000100001111,
    64'b0000000111000000000000000000100010000000010010000000000100001111,
    64'b0000000111000000000000000000010010000000010010000000001000001111,
    64'b0000000111000000000000000000010010000000010111111111101000001111,
    
    64'b1100000000000110000000000000000000000000000000000000000000000000,
    64'b1100000000000110000000000000000000000000000000000000000000000000,
    64'b1100000000000110000000000000000000000000000000000000000000000000,
    64'b1100000000000110000000000000000000000000000000000000000000000000,
    64'b1100000000000110000000000000000000000000000000000000000000000000,
    64'b1100000000000110000000000000000000000000000000000000000000000000,
    64'b1100000000000110000000000000000000000000000000000000000000000000,
    64'b1100000000000110000000000000000000000000000000000000000000000000,//7
    64'b1100000000000110000000000000000000000000000000000000000000000000,
    64'b1100000000000110000000000000000000000000000000000000000000000000,
    64'b1100000000000110000000000000000000000000000000000000000000000000,
    64'b1100000000000110000000000000000000000000000000000000000000000000,
    64'b1100000000000110000000000000000000000000000000000000000000000000,
    64'b1100000000000110000000000000000000000000000000000000000000000000,
    64'b1100000000000110000000000000000000000000000000000000000000000000,
    64'b1100000000000110000000000000000000000000000000000000000000000000,//7
    
    64'b0110000000001100000000000000010001110001110001000000010100001111,
    64'b0110000000001100000000000000010010001010001001000000010100001111,
    64'b0110000000001101100001100000100100000100000101000000010010001111,
    64'b0011000000011001010001010000100100000100000101000000010010001111,
    64'b0011000000011001001001001001000100000100000101000000010001000000,
    64'b0011000000011001000101000101000100000100000101000000010001000000,
    64'b0001100000110001000101000101000100000100000100100000100001000000,
    64'b0001100000110001001001001001000100000100000100100000100001000000,//7
    64'b0001100000110001010001010001000100000100000100100000100001000000,
    64'b0000110001100001100001100001000100000100000100100000100001000000,//9
    64'b0000110001100001000001000001000100000100000100010001000001000000,
    64'b0000110001100001000001000001000100000100000100010001000001000000,
    64'b0000011011000001000001000000100100000100000100010001000010001111,
    64'b0000011011000001000001000000100100000100000100001010000010001111,
    64'b0000001110000001000001000000010100000100000100000100000100001111,
    64'b0000000100000001000001000000010100000100000100000100000100001111
    };
    integer i;
    initial
     begin
      for(i=0;i<64;i=i+1)
        rom[i]=data[(4095-64*i)-:64];
     end
     
    assign F=rom[addr_Fre_Vopp];
 
    
endmodule
